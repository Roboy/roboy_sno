// darkroom.v

// Generated using ACDS version 17.1 590

`timescale 1 ps / 1 ps
module darkroom (
		input  wire       clk_clk,                           //                    clk.clk
		output wire       darkroom_0_conduit_end_mosi_o,     // darkroom_0_conduit_end.mosi_o
		output wire       darkroom_0_conduit_end_sck_o,      //                       .sck_o
		output wire       darkroom_0_conduit_end_ss_n_o,     //                       .ss_n_o
		input  wire       darkroom_0_conduit_end_trigger_me, //                       .trigger_me
		output wire [1:0] darkroom_0_conduit_end_sync_o,     //                       .sync_o
		inout  wire [1:0] darkroom_0_conduit_end_d_io,       //                       .d_io
		inout  wire [1:0] darkroom_0_conduit_end_e_io,       //                       .e_io
		input  wire       reset_reset_n                      //                  reset.reset_n
	);

	wire    rst_controller_reset_out_reset; // rst_controller:reset_out -> DarkRoom_0:reset_n

	DarkRoom #(
		.ENABLE_AVALON_INTERFACE (0),
		.ENABLE_SPI_TRANSMITTER  (1),
		.NUMBER_OF_SENSORS       (2),
		.CLK_SPEED               (32000000)
	) darkroom_0 (
		.reset_n     (~rst_controller_reset_out_reset),   //          reset.reset_n
		.mosi_o      (darkroom_0_conduit_end_mosi_o),     //    conduit_end.mosi_o
		.sck_o       (darkroom_0_conduit_end_sck_o),      //               .sck_o
		.ss_n_o      (darkroom_0_conduit_end_ss_n_o),     //               .ss_n_o
		.trigger_me  (darkroom_0_conduit_end_trigger_me), //               .trigger_me
		.sync_o      (darkroom_0_conduit_end_sync_o),     //               .sync_o
		.D_io        (darkroom_0_conduit_end_d_io),       //               .d_io
		.E_io        (darkroom_0_conduit_end_e_io),       //               .e_io
		.clock       (clk_clk),                           //     clock_sink.clk
		.address     (),                                  // avalon_slave_0.address
		.read        (),                                  //               .read
		.readdata    (),                                  //               .readdata
		.waitrequest ()                                   //               .waitrequest
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                 // reset_in0.reset
		.clk            (clk_clk),                        //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

endmodule
